constantVGA_inst : constantVGA PORT MAP (
		result	 => result_sig
	);
