BCD_Constant_inst : BCD_Constant PORT MAP (
		result	 => result_sig
	);
