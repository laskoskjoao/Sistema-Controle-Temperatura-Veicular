constant_ASCII_inst : constant_ASCII PORT MAP (
		result	 => result_sig
	);
