constControl_inst : constControl PORT MAP (
		result	 => result_sig
	);
