constante_teste_unidade_inst : constante_teste_unidade PORT MAP (
		result	 => result_sig
	);
