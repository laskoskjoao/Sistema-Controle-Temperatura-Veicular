constant_teste_dezena_inst : constant_teste_dezena PORT MAP (
		result	 => result_sig
	);
