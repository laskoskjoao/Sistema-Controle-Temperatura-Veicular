compare_inst : compare PORT MAP (
		dataa	 => dataa_sig,
		datab	 => datab_sig,
		aneb	 => aneb_sig
	);
