constante_teste_inst : constante_teste PORT MAP (
		result	 => result_sig
	);
