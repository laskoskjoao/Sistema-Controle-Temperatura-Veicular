compare_equal_inst : compare_equal PORT MAP (
		dataa	 => dataa_sig,
		datab	 => datab_sig,
		aeb	 => aeb_sig
	);
